`include "alu_if.sv"

package env_pkg; 
	`include "Packet.svh"
	`include "Scoreboard.svh"
	`include "monitor.svh"
	`include "driver.svh"
	`include "Stimulus_gen.svh"
endpackage 